`default_nettype none

module Not (
  output wire y,
  input wire a
);

  not(y, a);

endmodule


