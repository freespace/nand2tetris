`default_nettype none

module Not (
  output wire out,
  input wire a
);

  not(out, a);

endmodule


